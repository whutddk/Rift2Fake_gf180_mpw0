* NGSPICE file created from rift2Wrap.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

.subckt rift2Wrap io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0]
+ la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9]
+ la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15]
+ la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21]
+ la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28]
+ la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34]
+ la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40]
+ la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5]
+ la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8]
+ la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__519__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__338__A1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_363_ _048_ _134_ _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__329__A1 i_fake.lfsr_prng.io_out_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_294_ _082_ _083_ _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_346_ _056_ _117_ _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_277_ _055_ _056_ _059_ _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__532__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_200_ _141_ _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_329_ i_fake.lfsr_prng.io_out_15 i_fake.lfsr_prng.io_out_13 _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__527__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__347__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__374__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_84 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_73 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_62 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_95 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput20 net20 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput7 net7 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput31 net31 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput42 net42 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput53 net53 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_1_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__283__A1 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__535__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__C _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_362_ _023_ _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__329__A2 i_fake.lfsr_prng.io_out_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_293_ i_fake.lfsr_prng.io_out_0 _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__180__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__214__B _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__247__A1 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_345_ _068_ _122_ _123_ _119_ _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_276_ _071_ _058_ _063_ _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_328_ _110_ _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_259_ i_fake.lfsr_prng.io_out_4 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output12_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__312__B _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__358__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__268__I i_fake.lfsr_prng.io_out_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_74 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_63 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_85 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_96 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput10 net10 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput21 net21 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput8 net8 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput32 net32 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput43 net43 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput54 net54 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_1_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__178__I i_fake.lfsr_prng.io_out_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I la_oenb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__283__A2 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__387__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_361_ _033_ _129_ _133_ _132_ _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_292_ i_fake.lfsr_prng.io_out_1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_10_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__265__A2 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__320__B _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__247__A2 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_344_ _103_ _114_ _123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_275_ i_fake.lfsr_prng.io_out_7 _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__186__I i_fake.lfsr_prng.io_out_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_327_ _151_ _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_258_ i_fake.lfsr_prng.io_out_5 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_189_ i_fake.lfsr_prng.io_out_14 _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__359__A1 _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__307__C _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrift2Wrap_75 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_64 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_86 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_97 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput11 net11 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput9 net9 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput22 net22 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput33 net33 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput44 net44 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput55 net55 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__194__I i_fake.lfsr_prng.io_out_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_360_ _037_ _126_ _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_291_ _076_ _057_ _081_ _054_ net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__189__I i_fake.lfsr_prng.io_out_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__192__A2 _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_343_ _110_ _122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_274_ _057_ _059_ _064_ _070_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__377__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__292__I i_fake.lfsr_prng.io_out_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_326_ _104_ _084_ _109_ _054_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_257_ _048_ _028_ _053_ _054_ net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_188_ _143_ _147_ _152_ _155_ _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__310__A2 _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_309_ i_fake.lfsr_prng.io_out_3 _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__368__A2 _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__286__A1 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_65 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_76 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_87 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_98 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput12 net12 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput23 net23 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput34 net34 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput56 net56 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput45 net45 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__277__A1 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__201__A1 _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__295__I i_fake.lfsr_prng.io_out_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_290_ _066_ _067_ _062_ _072_ _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_342_ _098_ _111_ _121_ _119_ _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_273_ _066_ _067_ _069_ _169_ _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_325_ _093_ _094_ _089_ _099_ _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_256_ _019_ _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_187_ i_fake.lfsr_prng.io_out_14 _153_ _154_ _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__326__C _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_308_ _084_ _086_ _091_ _097_ net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_239_ _028_ _030_ _036_ _042_ net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__298__I i_fake.lfsr_prng.io_out_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output10_I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__210__A2 _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_66 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_77 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_88 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_99 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput13 net13 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 net24 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput57 net57 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_1_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput35 net35 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput46 net46 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__195__A1 i_fake.lfsr_prng.io_out_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I io_in[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_341_ _104_ _117_ _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_272_ _058_ _065_ _068_ _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_180 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__340__A1 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__322__A1 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_324_ _108_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_255_ _038_ _039_ _034_ _044_ _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_186_ i_fake.lfsr_prng.io_out_12 _154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__342__C _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_307_ _093_ _094_ _096_ _169_ _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_238_ _038_ _039_ _041_ _169_ _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrift2Wrap_78 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_89 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_67 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput14 net14 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput25 net25 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput58 net58 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput36 net36 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput47 net47 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__195__A2 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__345__C _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_340_ _088_ _111_ _120_ _119_ _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_27_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_271_ i_fake.lfsr_prng.io_out_4 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_170 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__322__A2 _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_323_ _024_ _107_ _108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_254_ _052_ net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_185_ i_fake.lfsr_prng.io_out_13 _153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__304__A2 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__231__A1 i_fake.lfsr_prng.io_out_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_306_ _085_ _092_ _095_ _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_237_ _029_ _037_ _040_ _041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_79 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_68 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput15 net15 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput37 net37 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput48 net48 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput26 net26 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput59 net59 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__361__C _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_270_ _060_ _061_ _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_160 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_171 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_537_ net24 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_322_ _103_ _084_ _090_ _094_ _093_ _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_253_ _024_ _051_ _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_7_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_184_ _151_ _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__231__A2 i_fake.lfsr_prng.io_out_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_305_ _083_ _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_236_ i_fake.lfsr_prng.io_out_8 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_144_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__380__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_219_ _023_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__364__C _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_69 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput38 net38 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput49 net49 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput16 net16 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput27 net27 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__361__A1 _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__359__C _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__352__A1 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output56_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_161 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_150 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_172 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_536_ net23 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__252__B1 _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_321_ _103_ _106_ _054_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_252_ _047_ _028_ _035_ _039_ _038_ _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_183_ _150_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_519_ net32 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__367__C _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_304_ _087_ _088_ _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_235_ _031_ _033_ _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__222__I i_fake.lfsr_prng.io_out_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_218_ _150_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput17 net17 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput28 net28 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput39 net39 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__198__A2 _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__370__A2 _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__352__A2 _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output9_I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__334__A2 _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_140 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_151 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_162 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_173 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_535_ net22 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__252__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__225__I i_fake.lfsr_prng.io_out_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_320_ _104_ _082_ _100_ _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_251_ _047_ _050_ _020_ net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_182_ _148_ net3 _149_ _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__234__A1 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_518_ net31 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__216__A1 _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_303_ _092_ _083_ _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_234_ _037_ i_fake.lfsr_prng.io_out_8 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_7_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_217_ _143_ _147_ _166_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__233__I i_fake.lfsr_prng.io_out_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__380__D _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput29 net29 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__375__D _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__228__I i_fake.lfsr_prng.io_out_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__511__I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__270__A2 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrift2Wrap_130 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_141 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_152 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_163 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_174 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_534_ net21 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_250_ _048_ _026_ _027_ _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_181_ net2 net3 _149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__234__A2 i_fake.lfsr_prng.io_out_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_517_ net30 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__383__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_379_ _005_ clknet_1_1__leaf_wb_clk_i i_fake.lfsr_prng.io_out_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__383__D _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__236__I i_fake.lfsr_prng.io_out_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_302_ i_fake.lfsr_prng.io_out_1 _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_233_ i_fake.lfsr_prng.io_out_9 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__378__D _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__373__A1 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_216_ _020_ _021_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__514__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput19 net19 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__355__A1 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__319__A1 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__386__D _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_120 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_142 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_131 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_153 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_164 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_175 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_533_ net20 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__522__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_180_ net1 _148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_516_ net29 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_378_ _004_ clknet_1_1__leaf_wb_clk_i i_fake.lfsr_prng.io_out_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__517__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_301_ _089_ _090_ _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_232_ _034_ _035_ _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__337__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__373__A2 _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_215_ _159_ _171_ _166_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__530__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__389__D _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__355__A2 _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__291__A1 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__346__A2 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__525__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_121 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_110 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_143 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_132 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_154 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_165 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_176 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_532_ net19 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output7_I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_515_ net28 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_377_ _003_ clknet_1_0__leaf_wb_clk_i i_fake.lfsr_prng.io_out_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__533__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__201__C _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_300_ i_fake.lfsr_prng.io_out_1 _083_ _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_231_ i_fake.lfsr_prng.io_out_9 i_fake.lfsr_prng.io_out_8 _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput1 io_in[28] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__528__I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__263__I i_fake.lfsr_prng.io_out_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_214_ _146_ _017_ _020_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__173__I i_fake.lfsr_prng.io_out_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__258__I i_fake.lfsr_prng.io_out_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__282__A2 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__386__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__536__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_100 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_111 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_144 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_133 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_122 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_155 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_166 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_177 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__271__I i_fake.lfsr_prng.io_out_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_531_ net18 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__182__A1 _148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__237__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_514_ net27 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__176__I i_fake.lfsr_prng.io_out_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_376_ _002_ clknet_1_0__leaf_wb_clk_i i_fake.lfsr_prng.io_out_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_230_ _031_ _033_ _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_359_ _026_ _129_ _131_ _132_ _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__300__A1 i_fake.lfsr_prng.io_out_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 la_data_in[0] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__367__A1 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_213_ _019_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrift2Wrap_101 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_112 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_145 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_134 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_123 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_156 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_167 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_178 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__191__A2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_530_ net17 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__182__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__237__A3 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__321__B _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__376__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output52_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_513_ net26 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_375_ _001_ clknet_1_0__leaf_wb_clk_i i_fake.lfsr_prng.io_out_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_358_ net4 _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_289_ _080_ net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__300__A2 _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 la_oenb[0] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__367__A2 _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_212_ net2 net3 _018_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__294__A1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__313__C _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__285__A1 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__249__A1 _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_102 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_135 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_124 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_113 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_146 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_157 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_168 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_179 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_512_ net25 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_374_ _000_ clknet_1_0__leaf_wb_clk_i i_fake.lfsr_prng.io_out_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output5_I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__293__I i_fake.lfsr_prng.io_out_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_357_ _027_ _126_ _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_288_ _024_ _079_ _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 wb_rst_i net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_211_ _148_ net3 _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__294__A2 _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__389__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__285__A2 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__249__A2 _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_103 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_136 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_125 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_114 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_158 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_147 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_169 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_144_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__330__A1 _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__321__A1 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_511_ net16 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_373_ _162_ _136_ _140_ _115_ _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__312__A1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__303__A1 _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_356_ _040_ _129_ _130_ _125_ _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_287_ _075_ _057_ _063_ _067_ _066_ _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_10_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_210_ _157_ _167_ _161_ _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_339_ _092_ _117_ _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__340__C _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__379__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_126 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_115 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_104 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_137 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_159 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_148 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_510_ net5 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_372_ _157_ _134_ _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__312__A2 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__303__A2 _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output50_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_355_ _075_ _114_ _130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_286_ _075_ _078_ _020_ net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__288__A1 _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__212__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_338_ _082_ _111_ _118_ _119_ _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_269_ _065_ i_fake.lfsr_prng.io_out_4 _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__338__C _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output13_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_127 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_116 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_105 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_138 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_149 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__330__A3 _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_371_ _145_ _136_ _139_ _115_ _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output43_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__230__A2 _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_354_ _110_ _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_285_ _076_ _055_ _056_ _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__212__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_337_ net4 _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_268_ i_fake.lfsr_prng.io_out_5 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_199_ _157_ _162_ _165_ _166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__360__A1 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__179__A1 _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__351__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_117 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_106 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_139 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_128 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__333__A1 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__306__A1 _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_370_ _153_ _134_ _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_353_ _071_ _122_ _128_ _125_ _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_284_ _061_ _063_ _077_ _062_ _070_ net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__302__I i_fake.lfsr_prng.io_out_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_336_ _100_ _117_ _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_267_ _062_ _063_ _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_198_ _141_ _142_ _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__188__B _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_319_ _088_ _090_ _105_ _089_ _097_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__360__A2 _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__179__A2 _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_107 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_118 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_129 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__333__A2 _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__286__B _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__260__A1 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__305__I _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__251__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__306__A2 _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__242__A1 _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__224__A1 _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__373__C _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_352_ _076_ _126_ _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_283_ _075_ _076_ _077_ _074_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__206__A1 _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__278__C _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_335_ _023_ _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_266_ i_fake.lfsr_prng.io_out_5 i_fake.lfsr_prng.io_out_4 _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_197_ _156_ _160_ _164_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__223__I i_fake.lfsr_prng.io_out_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_318_ _103_ _104_ _105_ _102_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_249_ _033_ _035_ _049_ _034_ _042_ net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output11_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__291__C _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_108 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_119 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output59_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__316__I _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I la_data_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__382__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_351_ _061_ _122_ _127_ _125_ _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_282_ _065_ _068_ _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_6_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__206__A2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_334_ _111_ _113_ _116_ _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_265_ _060_ _061_ _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_196_ _153_ _161_ _163_ _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__363__A1 _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_317_ _092_ _095_ _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__345__A1 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_248_ _047_ _048_ _049_ _046_ net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_179_ _145_ _146_ _147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__336__A1 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__381__D _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrift2Wrap_109 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__318__A1 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__376__D _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__512__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__332__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_350_ _065_ _126_ _127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_281_ _058_ _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__384__D _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_333_ _100_ _114_ _115_ _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_264_ i_fake.lfsr_prng.io_out_6 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__372__A2 _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_195_ i_fake.lfsr_prng.io_out_14 _162_ _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__363__A2 _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__520__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__379__D _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_316_ _085_ _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_247_ _037_ _040_ _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_178_ i_fake.lfsr_prng.io_out_15 _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__515__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__336__A2 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__335__I _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__318__A2 _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__387__D _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__209__A1 _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__523__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_280_ _060_ _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__518__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_332_ net4 _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_263_ i_fake.lfsr_prng.io_out_7 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_194_ i_fake.lfsr_prng.io_out_15 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_315_ _087_ _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_246_ _029_ _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_177_ _144_ _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__531__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_229_ _032_ _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__385__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__526__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__261__I i_fake.lfsr_prng.io_out_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__181__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output57_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__366__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__534__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_331_ _151_ _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_262_ i_fake.lfsr_prng.io_out_7 _058_ _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_193_ _142_ _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__348__A1 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_529_ net15 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__529__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__339__A1 _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__264__I i_fake.lfsr_prng.io_out_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_314_ _093_ _099_ _102_ _091_ net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_30_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__174__I i_fake.lfsr_prng.io_out_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_245_ _031_ _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_176_ i_fake.lfsr_prng.io_out_14 _144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__349__I _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__259__I i_fake.lfsr_prng.io_out_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__272__A3 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_228_ i_fake.lfsr_prng.io_out_10 _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__181__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__362__I _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__537__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__375__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__366__A2 _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_330_ _142_ _032_ _112_ _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__357__A2 _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_261_ i_fake.lfsr_prng.io_out_6 _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_192_ _157_ _146_ _159_ _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_528_ net14 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__284__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__339__A2 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_313_ _087_ _096_ _101_ _152_ _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_244_ _038_ _044_ _046_ _036_ net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_175_ _141_ _142_ _143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__266__A1 i_fake.lfsr_prng.io_out_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__257__A1 _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__275__I i_fake.lfsr_prng.io_out_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__248__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__185__I i_fake.lfsr_prng.io_out_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_227_ i_fake.lfsr_prng.io_out_11 _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__193__I _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_260_ _055_ _056_ _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_191_ _141_ _158_ _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_527_ net13 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_389_ _015_ clknet_1_0__leaf_wb_clk_i i_fake.lfsr_prng.io_out_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__388__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_312_ _082_ _100_ _086_ _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_14_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_243_ _031_ _041_ _045_ _152_ _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_174_ i_fake.lfsr_prng.io_out_12 _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__266__A2 i_fake.lfsr_prng.io_out_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__248__A2 _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_226_ i_fake.lfsr_prng.io_out_11 _029_ _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_209_ _145_ _165_ _016_ _156_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__320__A1 _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__369__A1 _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output55_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__333__B _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_190_ _154_ _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_526_ net12 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_388_ _014_ clknet_1_1__leaf_wb_clk_i i_fake.lfsr_prng.io_out_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_311_ i_fake.lfsr_prng.io_out_0 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_242_ _026_ _027_ _030_ _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_173_ i_fake.lfsr_prng.io_out_13 _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_225_ i_fake.lfsr_prng.io_out_10 _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__378__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__175__A2 _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__251__B _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_208_ _153_ _158_ _163_ _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__320__A2 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__297__I i_fake.lfsr_prng.io_out_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__369__A2 _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output48_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__296__A1 i_fake.lfsr_prng.io_out_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output8_I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__220__A1 _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__287__A1 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__211__A1 _148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__243__C _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_525_ net11 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_387_ _013_ clknet_1_1__leaf_wb_clk_i i_fake.lfsr_prng.io_out_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_310_ _098_ _085_ _090_ _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__238__C _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_241_ _043_ _029_ _035_ _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_224_ _026_ _027_ _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_207_ _170_ _172_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__296__A2 _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__211__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_524_ net10 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_386_ _012_ clknet_1_1__leaf_wb_clk_i i_fake.lfsr_prng.io_out_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__269__A2 i_fake.lfsr_prng.io_out_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_240_ i_fake.lfsr_prng.io_out_11 _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__187__A1 i_fake.lfsr_prng.io_out_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_369_ _167_ _136_ _138_ _115_ _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ i_fake.lfsr_prng.io_out_8 _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__341__A1 _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__323__A1 _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_206_ _145_ _158_ _171_ _172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__257__C _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output53_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_523_ net9 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_385_ _011_ clknet_1_0__leaf_wb_clk_i i_fake.lfsr_prng.io_out_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_368_ _161_ _134_ _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_299_ _087_ _088_ _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__350__A2 _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_222_ i_fake.lfsr_prng.io_out_9 _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__341__A2 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__323__A2 _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_205_ _146_ _167_ _171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__250__A1 _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__214__A1 _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__273__C _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__205__A1 _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_522_ net8 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_384_ _010_ clknet_1_1__leaf_wb_clk_i i_fake.lfsr_prng.io_out_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_90 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output6_I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_367_ _158_ _136_ _137_ _132_ _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_298_ i_fake.lfsr_prng.io_out_2 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__371__C _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_1__f_wb_clk_i clknet_0_wb_clk_i clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_221_ _163_ _022_ _025_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_204_ _143_ _166_ _170_ _164_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__311__I i_fake.lfsr_prng.io_out_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__250__A2 _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__232__A2 _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__299__A2 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__381__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__205__A2 _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_521_ net7 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_383_ _009_ clknet_1_1__leaf_wb_clk_i i_fake.lfsr_prng.io_out_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_80 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_91 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__371__A1 _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput60 net60 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__369__C _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_0__f_wb_clk_i clknet_0_wb_clk_i clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_366_ _047_ _114_ _137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_297_ i_fake.lfsr_prng.io_out_3 _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__344__A1 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_220_ _024_ _155_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__326__A1 _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__309__I i_fake.lfsr_prng.io_out_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__317__A1 _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_349_ _023_ _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__219__I _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__308__A1 _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_203_ _159_ _163_ _168_ _169_ _170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__241__A3 _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__374__D _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__227__I i_fake.lfsr_prng.io_out_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_520_ net6 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__199__A2 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_382_ _008_ clknet_1_0__leaf_wb_clk_i i_fake.lfsr_prng.io_out_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrift2Wrap_81 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_70 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_92 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__371__A2 _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput50 net50 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__510__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output51_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_365_ _110_ _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_296_ i_fake.lfsr_prng.io_out_3 _085_ _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__344__A2 _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__240__I i_fake.lfsr_prng.io_out_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__326__A2 _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__262__A1 i_fake.lfsr_prng.io_out_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_348_ _055_ _122_ _124_ _125_ _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_279_ _066_ _072_ _074_ _064_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_6_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__253__A1 _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__308__A2 _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__382__D _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_202_ _151_ _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__377__D _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__226__A1 i_fake.lfsr_prng.io_out_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__513__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_381_ _007_ clknet_1_1__leaf_wb_clk_i i_fake.lfsr_prng.io_out_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_82 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_71 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_93 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput5 net5 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput40 net40 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput51 net51 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__385__D _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_364_ _043_ _129_ _135_ _132_ _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_295_ i_fake.lfsr_prng.io_out_2 _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__521__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_347_ net4 _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_278_ _060_ _069_ _073_ _152_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__516__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__384__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_201_ _167_ _161_ _144_ _162_ _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__235__A2 _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__208__A2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__388__D _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__524__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_380_ _006_ clknet_1_1__leaf_wb_clk_i i_fake.lfsr_prng.io_out_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__356__A1 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_83 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_72 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xrift2Wrap_61 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrift2Wrap_94 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput6 net6 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput30 net30 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput52 net52 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput41 net41 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

